library IEEE;
use     IEEE.std_logic_1164.all;
use     IEEE.numeric_std.all;

entity FETCH is

  port (
    CLK         : in  std_logic;
    RST         : in  std_logic;
    PC_CURRENT  : in  std_logic_vector(31 downto 0);
    NOP         : in  std_logic;
    INSTRUCTION : out std_logic_vector(31 downto 0));
  
end entity FETCH;

architecture RTL of FETCH is
  
  signal S_MUX : std_logic_vector(31 downto 0);

  --  PROGRAMA 02:
  
  --1 MOV r0, #1
  -- "0000 00 1 1010 0 0000 0000 000001 000 000"  - CLK 4
  --2 MOV r1, #8
  -- "0000 00 1 1010 0 0001 0000 000001 000 011"  - CLK 5
  --3 SUB r2, r1, r0  
  -- "0000 00 0 0010 0 0010 0001 000000 000 000"  - CLK 6
  --4 STR M[10], r2
  -- "0000 01 1 00 1 0 0 0010 0000 000000001010"  - CLK 7
  --5 MOV LR, PC
  -- "0000 00 0 1010 0 1110 0000 001111 000 000"  - PC = 7;
  --6 NOP
  -- "0000 00 0 1010 0 0000 0000 000000 000 000"  - Besoin de NOP pour "prendre" le PC correct
  --7 CMP r2, #0
  -- "0000 00 1 1100 0 0000 0010 000000 000 000"  
  --8 BRANCH_EQ PC <- 12
  -- "0000 10 1 0 000000000000000000001100"       
  --9 SUBGT r2, r2, #1
  -- "1100 00 1 0010 1 0010 0010 000001 000 000"  
  --10 ADDLT r2, r2, #1
  -- "1011 00 1 0000 1 0010 0010 000001 000 000" 
  --11 MOV PC, LR
  -- "0000 00 0 1010 0 1111 0000 001110 000 000"  
  --12 LOAD M[10], r2
  -- "0000 01 1 00 0 0 0 0010 0000 000000001010"
  --13 MOV r2, r0, SLL#4
  -- "0000 00 0 1010 0 0010 0000 000000 000 100"
  --14 ADD r2, r2, r1
  -- "0000 00 0 0000 0 0010 0010 000001 000 000"
  --15 NOP
  -- "0000 00 0 1010 0 0000 0000 000000 000 000"
  --16 MOV LR, #1
  -- "0000 00 1 1010 0 1110 0000 000001 000 000"
  --17 MOV PC, LR
  -- "0000 00 0 1010 0 1111 0000 001110 000 000" 




  type TAB_ROM is array (0 to 63) of std_logic_vector(31 downto 0);
  constant MEM_INST : TAB_ROM :=
    (0  => "00000000000000000000000000000000", 1 => "00000011010000000000000001000000", 2 => "00000011010000010000000001000011",
     3  => "00000000010000100001000000000000", 4 => "00000110010000100000000000001010", 5 => "00000001010011100000001111000000",
     6  => "00000001010000000000000000000000", 7 => "00000011100000000010000000000000", 8 => "00001010000000000000000000001100",
     9  => "11000010010100100010000001000000", 10 => "10110010000100100010000001000000", 11 => "00000001010011110000001110000000",
     12 => "00000110000000100000000000001010", 13 => "00000001010000100000000000000100", 14 => "00000000000000100010000001000000",
     15 => "00000001010000000000000000000000", 16 => "00000011010011100000000001000000", 17 => "00000001010011110000001110000000",
     18 => "00000000000000000000000000000000", 19 => "00000000000000000000000000000000", 20 => "00000000000000000000000000000000",
     21 => "00000000000000000000000000000000", 22 => "00000000000000000000000000000000", 23 => "00000000000000000000000000000000",
     24 => "00000000000000000000000000000000", 25 => "00000000000000000000000000000000", 26 => "00000000000000000000000000000000",
     27 => "00000000000000000000000000000000", 28 => "00000000000000000000000000000000", 29 => "00000000000000000000000000000000",
     30 => "00000000000000000000000000000000", 31 => "00000000000000000000000000000000", 32 => "00000000000000000000000000000000",
     33 => "00000000000000000000000000000000", 34 => "00000000000000000000000000000000", 35 => "00000000000000000000000000000000",
     36 => "00000000000000000000000000000000", 37 => "00000000000000000000000000000000", 38 => "00000000000000000000000000000000",
     39 => "00000000000000000000000000000000", 40 => "00000000000000000000000000000000", 41 => "00000000000000000000000000000000",
     42 => "00000000000000000000000000000000", 43 => "00000000000000000000000000000000", 44 => "00000000000000000000000000000000",
     45 => "00000000000000000000000000000000", 46 => "00000000000000000000000000000000", 47 => "00000000000000000000000000000000",
     48 => "00000000000000000000000000000000", 49 => "00000000000000000000000000000000", 50 => "00000000000000000000000000000000",
     51 => "00000000000000000000000000000000", 52 => "00000000000000000000000000000000", 53 => "00000000000000000000000000000000",
     54 => "00000000000000000000000000000000", 55 => "00000000000000000000000000000000", 56 => "00000000000000000000000000000000",
     57 => "00000000000000000000000000000000", 58 => "00000000000000000000000000000000", 59 => "00000000000000000000000000000000",
     60 => "00000000000000000000000000000000", 61 => "00000000000000000000000000000000", 62 => "00000000000000000000000000000000",
     63 => "00000000000000000000000000000000");           
  
begin  -- architecture RTL

  -- MUX
  S_MUX <= MEM_INST(to_integer(unsigned(PC_CURRENT))) when NOP = '0' else
           "00000001010000000000000000000000";
 
  
  process (CLK, RST) is
  begin  -- process
    if CLK'event and CLK = '1' then  -- rising clock edge
      if RST = '1' then

        INSTRUCTION <= "00000000000000000000000000000000";

      else

        INSTRUCTION <= S_MUX;
        
      end if;
    end if;
  end process;
end architecture RTL;
